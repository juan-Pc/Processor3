--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:    00:10:46 10/17/2016 
-- Design Name:   
-- Module Name:   D:/Biblioteca/Documents/Procesador/Procesador32/MUXTB.vhd
-- Project Name:  Procesador
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: MUX
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY MUXTB IS
END MUXTB;
 
ARCHITECTURE behavior OF MUXTB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT MUX
    PORT(
         RfToMux : IN  std_logic_vector(31 downto 0);
         inm : IN  std_logic;
         seuToMux : IN  std_logic_vector(31 downto 0);
         MuxToAlu : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal RfToMux : std_logic_vector(31 downto 0) := (others => '0');
   signal inm : std_logic := '0';
   signal seuToMux : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal MuxToAlu : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MUX PORT MAP (
          RfToMux => RfToMux,
          inm => inm,
          seuToMux => seuToMux,
          MuxToAlu => MuxToAlu
        );

  

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      -- insert stimulus here 

      wait;
   end process;

END;
